* SPICE Model for LTK-0507-301-502 NPN Sensor

.subckt LTK0507 NPN_OUT VCC GND IN_LIGHT

* Sensor Parameters
.param V_ON = 10V   ; Min operating voltage
.param V_OFF = 30V  ; Max operating voltage
.param Imax = 100m  ; Max output current
.param Vdrop = 2V   ; Output voltage drop

* NPN Transistor Model (switching behavior)
Q1 NPN_OUT GND VCC NPNModel

* Light detection behavior (ON state when light is detected)
Vlight IN_LIGHT GND DC 0V ; Represents external light source
S1 NPN_OUT GND IN_LIGHT GND SW_LIGHT

.model NPNModel NPN(IS=1e-14 BF=100)

* Switching control based on light detection
.model SW_LIGHT SW(Ron=10m Roff=1Meg Vt=0.5V Vh=0.1V)

* Current Limitation for Output
R_limit NPN_OUT GND {Vdrop/Imax}

.ends LTK0507

* Simulation commands
* Example usage of the sensor model
X1 NPN_OUT VCC GND IN_LIGHT LTK0507

* Voltage sources
VCC VCC 0 DC 24V ; Power supply (between 10-30V)
VLIGHT IN_LIGHT 0 PULSE(0 1 0 1ms 1ms 2ms 4ms) ; Light source

* Simulation controls
.tran 0.1ms 10ms
.end
