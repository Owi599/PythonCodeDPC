*BSS138 N-Channel Logic Level Enhancement Mode Field Effect Transistor

.SUBCKT BSS138  D  G  S
* Pins: D - Drain, G - Gate, S - Source

* Model parameters
.PARAM Vth = 1.3V  ; Threshold voltage
.PARAM Kp = 0.12A/V^2  ; Transconductance parameter
.PARAM Lambda = 0.02V^-1  ; Channel length modulation
.PARAM Rd = 3.5Ohm  ; Drain resistance
.PARAM Rs = 3.5Ohm  ; Source resistance
.PARAM Cgd = 6pF  ; Gate-drain capacitance
.PARAM Cgs = 27pF  ; Gate-source capacitance
.PARAM Cds = 13pF  ; Drain-source capacitance

* MOSFET model
M1 D G S DMOS L=1u W=1u

.MODEL DMOS NMOS(Level=1, Vto={Vth}, Kp={Kp}, Lambda={Lambda})

* Resistors
Rd D drain {Rd}
Rs S source {Rs}

* Capacitors
Cgd G D {Cgd}
Cgs G S {Cgs}
Cds D S {Cds}

.ENDS BSS138